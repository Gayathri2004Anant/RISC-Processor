module my_and(
  input [31:0] in1,
  input [31:0] in2,
  output [31:0] out);
  
  and a0 (out[0], in1[0], in2[0]); 
  and a1 (out[1], in1[1], in2[1]); 
  and a2 (out[2], in1[2], in2[2]); 
  and a3 (out[3], in1[3], in2[3]); 
  and a4 (out[4], in1[4], in2[4]); 
  and a5 (out[5], in1[5], in2[5]); 
  and a6 (out[6], in1[6], in2[6]); 
  and a7 (out[7], in1[7], in2[7]); 
  and a8 (out[8], in1[8], in2[8]);
  and a9 (out[9], in1[9], in2[9]);
  and a10 (out[10], in1[10], in2[10]);
  and a11 (out[11], in1[11], in2[11]);
  and a12 (out[12], in1[12], in2[12]);
  and a13 (out[13], in1[13], in2[13]);
  and a14 (out[14], in1[14], in2[14]);
  and a15 (out[15], in1[15], in2[15]);
  and a16 (out[16], in1[16], in2[16]);
  and a17 (out[17], in1[17], in2[17]);
  and a18 (out[18], in1[18], in2[18]);
  and a19 (out[19], in1[19], in2[19]);
  and a20 (out[20], in1[20], in2[20]);
  and a21 (out[21], in1[21], in2[21]);
  and a22 (out[22], in1[22], in2[22]);
  and a23 (out[23], in1[23], in2[23]);
  and a24 (out[24], in1[24], in2[24]);
  and a25 (out[25], in1[25], in2[25]);
  and a26 (out[26], in1[26], in2[26]);
  and a27 (out[27], in1[27], in2[27]);
  and a28 (out[28], in1[28], in2[28]);
  and a29 (out[29], in1[29], in2[29]);
  and a30 (out[30], in1[30], in2[30]);
  and a31 (out[31], in1[31], in2[31]);
  
endmodule

module my_or(
  input [31:0] in1,
  input [31:0] in2,
  output [31:0] out);
  
  or a0 (out[0], in1[0], in2[0]); 
  or a1 (out[1], in1[1], in2[1]); 
  or a2 (out[2], in1[2], in2[2]); 
  or a3 (out[3], in1[3], in2[3]); 
  or a4 (out[4], in1[4], in2[4]); 
  or a5 (out[5], in1[5], in2[5]); 
  or a6 (out[6], in1[6], in2[6]); 
  or a7 (out[7], in1[7], in2[7]); 
  or a8 (out[8], in1[8], in2[8]);
  or a9 (out[9], in1[9], in2[9]);
  or a10 (out[10], in1[10], in2[10]);
  or a11 (out[11], in1[11], in2[11]);
  or a12 (out[12], in1[12], in2[12]);
  or a13 (out[13], in1[13], in2[13]);
  or a14 (out[14], in1[14], in2[14]);
  or a15 (out[15], in1[15], in2[15]);
  or a16 (out[16], in1[16], in2[16]);
  or a17 (out[17], in1[17], in2[17]);
  or a18 (out[18], in1[18], in2[18]);
  or a19 (out[19], in1[19], in2[19]);
  or a20 (out[20], in1[20], in2[20]);
  or a21 (out[21], in1[21], in2[21]);
  or a22 (out[22], in1[22], in2[22]);
  or a23 (out[23], in1[23], in2[23]);
  or a24 (out[24], in1[24], in2[24]);
  or a25 (out[25], in1[25], in2[25]);
  or a26 (out[26], in1[26], in2[26]);
  or a27 (out[27], in1[27], in2[27]);
  or a28 (out[28], in1[28], in2[28]);
  or a29 (out[29], in1[29], in2[29]);
  or a30 (out[30], in1[30], in2[30]);
  or a31 (out[31], in1[31], in2[31]);
  
endmodule

module my_xor(
  input [31:0] in1,
  input [31:0] in2,
  output [31:0] out);
  
  xor a0 (out[0], in1[0], in2[0]); 
  xor a1 (out[1], in1[1], in2[1]); 
  xor a2 (out[2], in1[2], in2[2]); 
  xor a3 (out[3], in1[3], in2[3]); 
  xor a4 (out[4], in1[4], in2[4]); 
  xor a5 (out[5], in1[5], in2[5]); 
  xor a6 (out[6], in1[6], in2[6]); 
  xor a7 (out[7], in1[7], in2[7]); 
  xor a8 (out[8], in1[8], in2[8]);
  xor a9 (out[9], in1[9], in2[9]);
  xor a10 (out[10], in1[10], in2[10]);
  xor a11 (out[11], in1[11], in2[11]);
  xor a12 (out[12], in1[12], in2[12]);
  xor a13 (out[13], in1[13], in2[13]);
  xor a14 (out[14], in1[14], in2[14]);
  xor a15 (out[15], in1[15], in2[15]);
  xor a16 (out[16], in1[16], in2[16]);
  xor a17 (out[17], in1[17], in2[17]);
  xor a18 (out[18], in1[18], in2[18]);
  xor a19 (out[19], in1[19], in2[19]);
  xor a20 (out[20], in1[20], in2[20]);
  xor a21 (out[21], in1[21], in2[21]);
  xor a22 (out[22], in1[22], in2[22]);
  xor a23 (out[23], in1[23], in2[23]);
  xor a24 (out[24], in1[24], in2[24]);
  xor a25 (out[25], in1[25], in2[25]);
  xor a26 (out[26], in1[26], in2[26]);
  xor a27 (out[27], in1[27], in2[27]);
  xor a28 (out[28], in1[28], in2[28]);
  xor a29 (out[29], in1[29], in2[29]);
  xor a30 (out[30], in1[30], in2[30]);
  xor a31 (out[31], in1[31], in2[31]);
  
endmodule

module my_not(
  input [31:0] in1,
  output [31:0] out);
  
  not a0 (out[0], in1[0]); 
  not a1 (out[1], in1[1]); 
  not a2 (out[2], in1[2]); 
  not a3 (out[3], in1[3]); 
  not a4 (out[4], in1[4]); 
  not a5 (out[5], in1[5]); 
  not a6 (out[6], in1[6]); 
  not a7 (out[7], in1[7]); 
  not a8 (out[8], in1[8]);
  not a9 (out[9], in1[9]);
  not a10 (out[10], in1[10]);
  not a11 (out[11], in1[11]);
  not a12 (out[12], in1[12]);
  not a13 (out[13], in1[13]);
  not a14 (out[14], in1[14]);
  not a15 (out[15], in1[15]);
  not a16 (out[16], in1[16]);
  not a17 (out[17], in1[17]);
  not a18 (out[18], in1[18]);
  not a19 (out[19], in1[19]);
  not a20 (out[20], in1[20]);
  not a21 (out[21], in1[21]);
  not a22 (out[22], in1[22]);
  not a23 (out[23], in1[23]);
  not a24 (out[24], in1[24]);
  not a25 (out[25], in1[25]);
  not a26 (out[26], in1[26]);
  not a27 (out[27], in1[27]);
  not a28 (out[28], in1[28]);
  not a29 (out[29], in1[29]);
  not a30 (out[30], in1[30]);
  not a31 (out[31], in1[31]);
  
endmodule

module my_nor(
  input [31:0] in1,
  input [31:0] in2,
  output [31:0] out);

wire [31:0] temp;
my_or o (in1, in2, temp);
my_not n (temp, out);

endmodule