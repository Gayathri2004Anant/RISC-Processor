module right_shift_arith(input [31:0] in1, input [31:0] in2, output [31:0] out);
        wire [32:0] temp0;
		wire [32:0] temp1;
		wire [32:0] temp2;
		wire [32:0] temp3;
		wire [32:0] temp4;
		wire [32:0] temp5;
		wire [32:0] temp6;
		wire [32:0] temp7;
		wire [32:0] temp8;
		wire [32:0] temp9;
		wire [32:0] temp10;
		wire [32:0] temp11;
		wire [32:0] temp12;
		wire [32:0] temp13;
		wire [32:0] temp14;
		wire [32:0] temp15;
		wire [32:0] temp16;
		wire [32:0] temp17;
		wire [32:0] temp18;
		wire [32:0] temp19;
		wire [32:0] temp20;
		wire [32:0] temp21;
		wire [32:0] temp22;
		wire [32:0] temp23;
		wire [32:0] temp24;
		wire [32:0] temp25;
		wire [32:0] temp26;
		wire [32:0] temp27;
		wire [32:0] temp28;
		wire [32:0] temp29;
		wire [32:0] temp30;
		wire [32:0] temp31;
		assign temp0 = in1;

		assign temp1[31] = in1[31];
		assign temp1[30:0] = in1[31:1];
		
		assign temp2[29:0] = in1[31:2];
assign temp2[31] = in1[31];
assign temp2[30] = in1[31];
assign temp3[28:0] = in1[31:3];
assign temp3[31] = in1[31];
assign temp3[30] = in1[31];
assign temp3[29] = in1[31];
assign temp4[27:0] = in1[31:4];
assign temp4[31] = in1[31];
assign temp4[30] = in1[31];
assign temp4[29] = in1[31];
assign temp4[28] = in1[31];
assign temp5[26:0] = in1[31:5];
assign temp5[31] = in1[31];
assign temp5[30] = in1[31];
assign temp5[29] = in1[31];
assign temp5[28] = in1[31];
assign temp5[27] = in1[31];
assign temp6[25:0] = in1[31:6];
assign temp6[31] = in1[31];
assign temp6[30] = in1[31];
assign temp6[29] = in1[31];
assign temp6[28] = in1[31];
assign temp6[27] = in1[31];
assign temp6[26] = in1[31];
assign temp7[24:0] = in1[31:7];
assign temp7[31] = in1[31];
assign temp7[30] = in1[31];
assign temp7[29] = in1[31];
assign temp7[28] = in1[31];
assign temp7[27] = in1[31];
assign temp7[26] = in1[31];
assign temp7[25] = in1[31];
assign temp8[23:0] = in1[31:8];
assign temp8[31] = in1[31];
assign temp8[30] = in1[31];
assign temp8[29] = in1[31];
assign temp8[28] = in1[31];
assign temp8[27] = in1[31];
assign temp8[26] = in1[31];
assign temp8[25] = in1[31];
assign temp8[24] = in1[31];
assign temp9[22:0] = in1[31:9];
assign temp9[31] = in1[31];
assign temp9[30] = in1[31];
assign temp9[29] = in1[31];
assign temp9[28] = in1[31];
assign temp9[27] = in1[31];
assign temp9[26] = in1[31];
assign temp9[25] = in1[31];
assign temp9[24] = in1[31];
assign temp9[23] = in1[31];
assign temp10[21:0] = in1[31:10];
assign temp10[31] = in1[31];
assign temp10[30] = in1[31];
assign temp10[29] = in1[31];
assign temp10[28] = in1[31];
assign temp10[27] = in1[31];
assign temp10[26] = in1[31];
assign temp10[25] = in1[31];
assign temp10[24] = in1[31];
assign temp10[23] = in1[31];
assign temp10[22] = in1[31];
assign temp11[20:0] = in1[31:11];
assign temp11[31] = in1[31];
assign temp11[30] = in1[31];
assign temp11[29] = in1[31];
assign temp11[28] = in1[31];
assign temp11[27] = in1[31];
assign temp11[26] = in1[31];
assign temp11[25] = in1[31];
assign temp11[24] = in1[31];
assign temp11[23] = in1[31];
assign temp11[22] = in1[31];
assign temp11[21] = in1[31];
assign temp12[19:0] = in1[31:12];
assign temp12[31] = in1[31];
assign temp12[30] = in1[31];
assign temp12[29] = in1[31];
assign temp12[28] = in1[31];
assign temp12[27] = in1[31];
assign temp12[26] = in1[31];
assign temp12[25] = in1[31];
assign temp12[24] = in1[31];
assign temp12[23] = in1[31];
assign temp12[22] = in1[31];
assign temp12[21] = in1[31];
assign temp12[20] = in1[31];
assign temp13[18:0] = in1[31:13];
assign temp13[31] = in1[31];
assign temp13[30] = in1[31];
assign temp13[29] = in1[31];
assign temp13[28] = in1[31];
assign temp13[27] = in1[31];
assign temp13[26] = in1[31];
assign temp13[25] = in1[31];
assign temp13[24] = in1[31];
assign temp13[23] = in1[31];
assign temp13[22] = in1[31];
assign temp13[21] = in1[31];
assign temp13[20] = in1[31];
assign temp13[19] = in1[31];
assign temp14[17:0] = in1[31:14];
assign temp14[31] = in1[31];
assign temp14[30] = in1[31];
assign temp14[29] = in1[31];
assign temp14[28] = in1[31];
assign temp14[27] = in1[31];
assign temp14[26] = in1[31];
assign temp14[25] = in1[31];
assign temp14[24] = in1[31];
assign temp14[23] = in1[31];
assign temp14[22] = in1[31];
assign temp14[21] = in1[31];
assign temp14[20] = in1[31];
assign temp14[19] = in1[31];
assign temp14[18] = in1[31];
assign temp15[16:0] = in1[31:15];
assign temp15[31] = in1[31];
assign temp15[30] = in1[31];
assign temp15[29] = in1[31];
assign temp15[28] = in1[31];
assign temp15[27] = in1[31];
assign temp15[26] = in1[31];
assign temp15[25] = in1[31];
assign temp15[24] = in1[31];
assign temp15[23] = in1[31];
assign temp15[22] = in1[31];
assign temp15[21] = in1[31];
assign temp15[20] = in1[31];
assign temp15[19] = in1[31];
assign temp15[18] = in1[31];
assign temp15[17] = in1[31];
assign temp16[15:0] = in1[31:16];
assign temp16[31] = in1[31];
assign temp16[30] = in1[31];
assign temp16[29] = in1[31];
assign temp16[28] = in1[31];
assign temp16[27] = in1[31];
assign temp16[26] = in1[31];
assign temp16[25] = in1[31];
assign temp16[24] = in1[31];
assign temp16[23] = in1[31];
assign temp16[22] = in1[31];
assign temp16[21] = in1[31];
assign temp16[20] = in1[31];
assign temp16[19] = in1[31];
assign temp16[18] = in1[31];
assign temp16[17] = in1[31];
assign temp16[16] = in1[31];
assign temp17[14:0] = in1[31:17];
assign temp17[31] = in1[31];
assign temp17[30] = in1[31];
assign temp17[29] = in1[31];
assign temp17[28] = in1[31];
assign temp17[27] = in1[31];
assign temp17[26] = in1[31];
assign temp17[25] = in1[31];
assign temp17[24] = in1[31];
assign temp17[23] = in1[31];
assign temp17[22] = in1[31];
assign temp17[21] = in1[31];
assign temp17[20] = in1[31];
assign temp17[19] = in1[31];
assign temp17[18] = in1[31];
assign temp17[17] = in1[31];
assign temp17[16] = in1[31];
assign temp17[15] = in1[31];
assign temp18[13:0] = in1[31:18];
assign temp18[31] = in1[31];
assign temp18[30] = in1[31];
assign temp18[29] = in1[31];
assign temp18[28] = in1[31];
assign temp18[27] = in1[31];
assign temp18[26] = in1[31];
assign temp18[25] = in1[31];
assign temp18[24] = in1[31];
assign temp18[23] = in1[31];
assign temp18[22] = in1[31];
assign temp18[21] = in1[31];
assign temp18[20] = in1[31];
assign temp18[19] = in1[31];
assign temp18[18] = in1[31];
assign temp18[17] = in1[31];
assign temp18[16] = in1[31];
assign temp18[15] = in1[31];
assign temp18[14] = in1[31];
assign temp19[12:0] = in1[31:19];
assign temp19[31] = in1[31];
assign temp19[30] = in1[31];
assign temp19[29] = in1[31];
assign temp19[28] = in1[31];
assign temp19[27] = in1[31];
assign temp19[26] = in1[31];
assign temp19[25] = in1[31];
assign temp19[24] = in1[31];
assign temp19[23] = in1[31];
assign temp19[22] = in1[31];
assign temp19[21] = in1[31];
assign temp19[20] = in1[31];
assign temp19[19] = in1[31];
assign temp19[18] = in1[31];
assign temp19[17] = in1[31];
assign temp19[16] = in1[31];
assign temp19[15] = in1[31];
assign temp19[14] = in1[31];
assign temp19[13] = in1[31];
assign temp20[11:0] = in1[31:20];
assign temp20[31] = in1[31];
assign temp20[30] = in1[31];
assign temp20[29] = in1[31];
assign temp20[28] = in1[31];
assign temp20[27] = in1[31];
assign temp20[26] = in1[31];
assign temp20[25] = in1[31];
assign temp20[24] = in1[31];
assign temp20[23] = in1[31];
assign temp20[22] = in1[31];
assign temp20[21] = in1[31];
assign temp20[20] = in1[31];
assign temp20[19] = in1[31];
assign temp20[18] = in1[31];
assign temp20[17] = in1[31];
assign temp20[16] = in1[31];
assign temp20[15] = in1[31];
assign temp20[14] = in1[31];
assign temp20[13] = in1[31];
assign temp20[12] = in1[31];
assign temp21[10:0] = in1[31:21];
assign temp21[31] = in1[31];
assign temp21[30] = in1[31];
assign temp21[29] = in1[31];
assign temp21[28] = in1[31];
assign temp21[27] = in1[31];
assign temp21[26] = in1[31];
assign temp21[25] = in1[31];
assign temp21[24] = in1[31];
assign temp21[23] = in1[31];
assign temp21[22] = in1[31];
assign temp21[21] = in1[31];
assign temp21[20] = in1[31];
assign temp21[19] = in1[31];
assign temp21[18] = in1[31];
assign temp21[17] = in1[31];
assign temp21[16] = in1[31];
assign temp21[15] = in1[31];
assign temp21[14] = in1[31];
assign temp21[13] = in1[31];
assign temp21[12] = in1[31];
assign temp21[11] = in1[31];
assign temp22[9:0] = in1[31:22];
assign temp22[31] = in1[31];
assign temp22[30] = in1[31];
assign temp22[29] = in1[31];
assign temp22[28] = in1[31];
assign temp22[27] = in1[31];
assign temp22[26] = in1[31];
assign temp22[25] = in1[31];
assign temp22[24] = in1[31];
assign temp22[23] = in1[31];
assign temp22[22] = in1[31];
assign temp22[21] = in1[31];
assign temp22[20] = in1[31];
assign temp22[19] = in1[31];
assign temp22[18] = in1[31];
assign temp22[17] = in1[31];
assign temp22[16] = in1[31];
assign temp22[15] = in1[31];
assign temp22[14] = in1[31];
assign temp22[13] = in1[31];
assign temp22[12] = in1[31];
assign temp22[11] = in1[31];
assign temp22[10] = in1[31];
assign temp23[8:0] = in1[31:23];
assign temp23[31] = in1[31];
assign temp23[30] = in1[31];
assign temp23[29] = in1[31];
assign temp23[28] = in1[31];
assign temp23[27] = in1[31];
assign temp23[26] = in1[31];
assign temp23[25] = in1[31];
assign temp23[24] = in1[31];
assign temp23[23] = in1[31];
assign temp23[22] = in1[31];
assign temp23[21] = in1[31];
assign temp23[20] = in1[31];
assign temp23[19] = in1[31];
assign temp23[18] = in1[31];
assign temp23[17] = in1[31];
assign temp23[16] = in1[31];
assign temp23[15] = in1[31];
assign temp23[14] = in1[31];
assign temp23[13] = in1[31];
assign temp23[12] = in1[31];
assign temp23[11] = in1[31];
assign temp23[10] = in1[31];
assign temp23[9] = in1[31];
assign temp24[7:0] = in1[31:24];
assign temp24[31] = in1[31];
assign temp24[30] = in1[31];
assign temp24[29] = in1[31];
assign temp24[28] = in1[31];
assign temp24[27] = in1[31];
assign temp24[26] = in1[31];
assign temp24[25] = in1[31];
assign temp24[24] = in1[31];
assign temp24[23] = in1[31];
assign temp24[22] = in1[31];
assign temp24[21] = in1[31];
assign temp24[20] = in1[31];
assign temp24[19] = in1[31];
assign temp24[18] = in1[31];
assign temp24[17] = in1[31];
assign temp24[16] = in1[31];
assign temp24[15] = in1[31];
assign temp24[14] = in1[31];
assign temp24[13] = in1[31];
assign temp24[12] = in1[31];
assign temp24[11] = in1[31];
assign temp24[10] = in1[31];
assign temp24[9] = in1[31];
assign temp24[8] = in1[31];
assign temp25[6:0] = in1[31:25];
assign temp25[31] = in1[31];
assign temp25[30] = in1[31];
assign temp25[29] = in1[31];
assign temp25[28] = in1[31];
assign temp25[27] = in1[31];
assign temp25[26] = in1[31];
assign temp25[25] = in1[31];
assign temp25[24] = in1[31];
assign temp25[23] = in1[31];
assign temp25[22] = in1[31];
assign temp25[21] = in1[31];
assign temp25[20] = in1[31];
assign temp25[19] = in1[31];
assign temp25[18] = in1[31];
assign temp25[17] = in1[31];
assign temp25[16] = in1[31];
assign temp25[15] = in1[31];
assign temp25[14] = in1[31];
assign temp25[13] = in1[31];
assign temp25[12] = in1[31];
assign temp25[11] = in1[31];
assign temp25[10] = in1[31];
assign temp25[9] = in1[31];
assign temp25[8] = in1[31];
assign temp25[7] = in1[31];
assign temp26[5:0] = in1[31:26];
assign temp26[31] = in1[31];
assign temp26[30] = in1[31];
assign temp26[29] = in1[31];
assign temp26[28] = in1[31];
assign temp26[27] = in1[31];
assign temp26[26] = in1[31];
assign temp26[25] = in1[31];
assign temp26[24] = in1[31];
assign temp26[23] = in1[31];
assign temp26[22] = in1[31];
assign temp26[21] = in1[31];
assign temp26[20] = in1[31];
assign temp26[19] = in1[31];
assign temp26[18] = in1[31];
assign temp26[17] = in1[31];
assign temp26[16] = in1[31];
assign temp26[15] = in1[31];
assign temp26[14] = in1[31];
assign temp26[13] = in1[31];
assign temp26[12] = in1[31];
assign temp26[11] = in1[31];
assign temp26[10] = in1[31];
assign temp26[9] = in1[31];
assign temp26[8] = in1[31];
assign temp26[7] = in1[31];
assign temp26[6] = in1[31];
assign temp27[4:0] = in1[31:27];
assign temp27[31] = in1[31];
assign temp27[30] = in1[31];
assign temp27[29] = in1[31];
assign temp27[28] = in1[31];
assign temp27[27] = in1[31];
assign temp27[26] = in1[31];
assign temp27[25] = in1[31];
assign temp27[24] = in1[31];
assign temp27[23] = in1[31];
assign temp27[22] = in1[31];
assign temp27[21] = in1[31];
assign temp27[20] = in1[31];
assign temp27[19] = in1[31];
assign temp27[18] = in1[31];
assign temp27[17] = in1[31];
assign temp27[16] = in1[31];
assign temp27[15] = in1[31];
assign temp27[14] = in1[31];
assign temp27[13] = in1[31];
assign temp27[12] = in1[31];
assign temp27[11] = in1[31];
assign temp27[10] = in1[31];
assign temp27[9] = in1[31];
assign temp27[8] = in1[31];
assign temp27[7] = in1[31];
assign temp27[6] = in1[31];
assign temp27[5] = in1[31];
assign temp28[3:0] = in1[31:28];
assign temp28[31] = in1[31];
assign temp28[30] = in1[31];
assign temp28[29] = in1[31];
assign temp28[28] = in1[31];
assign temp28[27] = in1[31];
assign temp28[26] = in1[31];
assign temp28[25] = in1[31];
assign temp28[24] = in1[31];
assign temp28[23] = in1[31];
assign temp28[22] = in1[31];
assign temp28[21] = in1[31];
assign temp28[20] = in1[31];
assign temp28[19] = in1[31];
assign temp28[18] = in1[31];
assign temp28[17] = in1[31];
assign temp28[16] = in1[31];
assign temp28[15] = in1[31];
assign temp28[14] = in1[31];
assign temp28[13] = in1[31];
assign temp28[12] = in1[31];
assign temp28[11] = in1[31];
assign temp28[10] = in1[31];
assign temp28[9] = in1[31];
assign temp28[8] = in1[31];
assign temp28[7] = in1[31];
assign temp28[6] = in1[31];
assign temp28[5] = in1[31];
assign temp28[4] = in1[31];
assign temp29[2:0] = in1[31:29];
assign temp29[31] = in1[31];
assign temp29[30] = in1[31];
assign temp29[29] = in1[31];
assign temp29[28] = in1[31];
assign temp29[27] = in1[31];
assign temp29[26] = in1[31];
assign temp29[25] = in1[31];
assign temp29[24] = in1[31];
assign temp29[23] = in1[31];
assign temp29[22] = in1[31];
assign temp29[21] = in1[31];
assign temp29[20] = in1[31];
assign temp29[19] = in1[31];
assign temp29[18] = in1[31];
assign temp29[17] = in1[31];
assign temp29[16] = in1[31];
assign temp29[15] = in1[31];
assign temp29[14] = in1[31];
assign temp29[13] = in1[31];
assign temp29[12] = in1[31];
assign temp29[11] = in1[31];
assign temp29[10] = in1[31];
assign temp29[9] = in1[31];
assign temp29[8] = in1[31];
assign temp29[7] = in1[31];
assign temp29[6] = in1[31];
assign temp29[5] = in1[31];
assign temp29[4] = in1[31];
assign temp29[3] = in1[31];
assign temp30[1:0] = in1[31:30];
assign temp30[31] = in1[31];
assign temp30[30] = in1[31];
assign temp30[29] = in1[31];
assign temp30[28] = in1[31];
assign temp30[27] = in1[31];
assign temp30[26] = in1[31];
assign temp30[25] = in1[31];
assign temp30[24] = in1[31];
assign temp30[23] = in1[31];
assign temp30[22] = in1[31];
assign temp30[21] = in1[31];
assign temp30[20] = in1[31];
assign temp30[19] = in1[31];
assign temp30[18] = in1[31];
assign temp30[17] = in1[31];
assign temp30[16] = in1[31];
assign temp30[15] = in1[31];
assign temp30[14] = in1[31];
assign temp30[13] = in1[31];
assign temp30[12] = in1[31];
assign temp30[11] = in1[31];
assign temp30[10] = in1[31];
assign temp30[9] = in1[31];
assign temp30[8] = in1[31];
assign temp30[7] = in1[31];
assign temp30[6] = in1[31];
assign temp30[5] = in1[31];
assign temp30[4] = in1[31];
assign temp30[3] = in1[31];
assign temp30[2] = in1[31];
assign temp31[0:0] = in1[31:31];
assign temp31[31] = in1[31];
assign temp31[30] = in1[31];
assign temp31[29] = in1[31];
assign temp31[28] = in1[31];
assign temp31[27] = in1[31];
assign temp31[26] = in1[31];
assign temp31[25] = in1[31];
assign temp31[24] = in1[31];
assign temp31[23] = in1[31];
assign temp31[22] = in1[31];
assign temp31[21] = in1[31];
assign temp31[20] = in1[31];
assign temp31[19] = in1[31];
assign temp31[18] = in1[31];
assign temp31[17] = in1[31];
assign temp31[16] = in1[31];
assign temp31[15] = in1[31];
assign temp31[14] = in1[31];
assign temp31[13] = in1[31];
assign temp31[12] = in1[31];
assign temp31[11] = in1[31];
assign temp31[10] = in1[31];
assign temp31[9] = in1[31];
assign temp31[8] = in1[31];
assign temp31[7] = in1[31];
assign temp31[6] = in1[31];
assign temp31[5] = in1[31];
assign temp31[4] = in1[31];
assign temp31[3] = in1[31];
assign temp31[2] = in1[31];
assign temp31[1] = in1[31];


			 
	 mux32to1 m0({temp31[0], temp30[0], temp29[0], temp28[0], temp27[0], temp26[0], temp25[0], temp24[0], temp23[0], temp22[0], temp21[0], temp20[0], temp19[0], temp18[0], temp17[0], temp16[0], temp15[0], temp14[0], temp13[0], temp12[0], temp11[0], temp10[0], temp9[0], temp8[0], temp7[0], temp6[0], temp5[0], temp4[0], temp3[0], temp2[0], temp1[0], temp0[0]}, in2[4:0], out[0]);
mux32to1 m1({temp31[1], temp30[1], temp29[1], temp28[1], temp27[1], temp26[1], temp25[1], temp24[1], temp23[1], temp22[1], temp21[1], temp20[1], temp19[1], temp18[1], temp17[1], temp16[1], temp15[1], temp14[1], temp13[1], temp12[1], temp11[1], temp10[1], temp9[1], temp8[1], temp7[1], temp6[1], temp5[1], temp4[1], temp3[1], temp2[1], temp1[1], temp0[1]}, in2[4:0], out[1]);
mux32to1 m2({temp31[2], temp30[2], temp29[2], temp28[2], temp27[2], temp26[2], temp25[2], temp24[2], temp23[2], temp22[2], temp21[2], temp20[2], temp19[2], temp18[2], temp17[2], temp16[2], temp15[2], temp14[2], temp13[2], temp12[2], temp11[2], temp10[2], temp9[2], temp8[2], temp7[2], temp6[2], temp5[2], temp4[2], temp3[2], temp2[2], temp1[2], temp0[2]}, in2[4:0], out[2]);
mux32to1 m3({temp31[3], temp30[3], temp29[3], temp28[3], temp27[3], temp26[3], temp25[3], temp24[3], temp23[3], temp22[3], temp21[3], temp20[3], temp19[3], temp18[3], temp17[3], temp16[3], temp15[3], temp14[3], temp13[3], temp12[3], temp11[3], temp10[3], temp9[3], temp8[3], temp7[3], temp6[3], temp5[3], temp4[3], temp3[3], temp2[3], temp1[3], temp0[3]}, in2[4:0], out[3]);
mux32to1 m4({temp31[4], temp30[4], temp29[4], temp28[4], temp27[4], temp26[4], temp25[4], temp24[4], temp23[4], temp22[4], temp21[4], temp20[4], temp19[4], temp18[4], temp17[4], temp16[4], temp15[4], temp14[4], temp13[4], temp12[4], temp11[4], temp10[4], temp9[4], temp8[4], temp7[4], temp6[4], temp5[4], temp4[4], temp3[4], temp2[4], temp1[4], temp0[4]}, in2[4:0], out[4]);
mux32to1 m5({temp31[5], temp30[5], temp29[5], temp28[5], temp27[5], temp26[5], temp25[5], temp24[5], temp23[5], temp22[5], temp21[5], temp20[5], temp19[5], temp18[5], temp17[5], temp16[5], temp15[5], temp14[5], temp13[5], temp12[5], temp11[5], temp10[5], temp9[5], temp8[5], temp7[5], temp6[5], temp5[5], temp4[5], temp3[5], temp2[5], temp1[5], temp0[5]}, in2[4:0], out[5]);
mux32to1 m6({temp31[6], temp30[6], temp29[6], temp28[6], temp27[6], temp26[6], temp25[6], temp24[6], temp23[6], temp22[6], temp21[6], temp20[6], temp19[6], temp18[6], temp17[6], temp16[6], temp15[6], temp14[6], temp13[6], temp12[6], temp11[6], temp10[6], temp9[6], temp8[6], temp7[6], temp6[6], temp5[6], temp4[6], temp3[6], temp2[6], temp1[6], temp0[6]}, in2[4:0], out[6]);
mux32to1 m7({temp31[7], temp30[7], temp29[7], temp28[7], temp27[7], temp26[7], temp25[7], temp24[7], temp23[7], temp22[7], temp21[7], temp20[7], temp19[7], temp18[7], temp17[7], temp16[7], temp15[7], temp14[7], temp13[7], temp12[7], temp11[7], temp10[7], temp9[7], temp8[7], temp7[7], temp6[7], temp5[7], temp4[7], temp3[7], temp2[7], temp1[7], temp0[7]}, in2[4:0], out[7]);
mux32to1 m8({temp31[8], temp30[8], temp29[8], temp28[8], temp27[8], temp26[8], temp25[8], temp24[8], temp23[8], temp22[8], temp21[8], temp20[8], temp19[8], temp18[8], temp17[8], temp16[8], temp15[8], temp14[8], temp13[8], temp12[8], temp11[8], temp10[8], temp9[8], temp8[8], temp7[8], temp6[8], temp5[8], temp4[8], temp3[8], temp2[8], temp1[8], temp0[8]}, in2[4:0], out[8]);
mux32to1 m9({temp31[9], temp30[9], temp29[9], temp28[9], temp27[9], temp26[9], temp25[9], temp24[9], temp23[9], temp22[9], temp21[9], temp20[9], temp19[9], temp18[9], temp17[9], temp16[9], temp15[9], temp14[9], temp13[9], temp12[9], temp11[9], temp10[9], temp9[9], temp8[9], temp7[9], temp6[9], temp5[9], temp4[9], temp3[9], temp2[9], temp1[9], temp0[9]}, in2[4:0], out[9]);
mux32to1 m10({temp31[10], temp30[10], temp29[10], temp28[10], temp27[10], temp26[10], temp25[10], temp24[10], temp23[10], temp22[10], temp21[10], temp20[10], temp19[10], temp18[10], temp17[10], temp16[10], temp15[10], temp14[10], temp13[10], temp12[10], temp11[10], temp10[10], temp9[10], temp8[10], temp7[10], temp6[10], temp5[10], temp4[10], temp3[10], temp2[10], temp1[10], temp0[10]}, in2[4:0], out[10]);
mux32to1 m11({temp31[11], temp30[11], temp29[11], temp28[11], temp27[11], temp26[11], temp25[11], temp24[11], temp23[11], temp22[11], temp21[11], temp20[11], temp19[11], temp18[11], temp17[11], temp16[11], temp15[11], temp14[11], temp13[11], temp12[11], temp11[11], temp10[11], temp9[11], temp8[11], temp7[11], temp6[11], temp5[11], temp4[11], temp3[11], temp2[11], temp1[11], temp0[11]}, in2[4:0], out[11]);
mux32to1 m12({temp31[12], temp30[12], temp29[12], temp28[12], temp27[12], temp26[12], temp25[12], temp24[12], temp23[12], temp22[12], temp21[12], temp20[12], temp19[12], temp18[12], temp17[12], temp16[12], temp15[12], temp14[12], temp13[12], temp12[12], temp11[12], temp10[12], temp9[12], temp8[12], temp7[12], temp6[12], temp5[12], temp4[12], temp3[12], temp2[12], temp1[12], temp0[12]}, in2[4:0], out[12]);
mux32to1 m13({temp31[13], temp30[13], temp29[13], temp28[13], temp27[13], temp26[13], temp25[13], temp24[13], temp23[13], temp22[13], temp21[13], temp20[13], temp19[13], temp18[13], temp17[13], temp16[13], temp15[13], temp14[13], temp13[13], temp12[13], temp11[13], temp10[13], temp9[13], temp8[13], temp7[13], temp6[13], temp5[13], temp4[13], temp3[13], temp2[13], temp1[13], temp0[13]}, in2[4:0], out[13]);
mux32to1 m14({temp31[14], temp30[14], temp29[14], temp28[14], temp27[14], temp26[14], temp25[14], temp24[14], temp23[14], temp22[14], temp21[14], temp20[14], temp19[14], temp18[14], temp17[14], temp16[14], temp15[14], temp14[14], temp13[14], temp12[14], temp11[14], temp10[14], temp9[14], temp8[14], temp7[14], temp6[14], temp5[14], temp4[14], temp3[14], temp2[14], temp1[14], temp0[14]}, in2[4:0], out[14]);
mux32to1 m15({temp31[15], temp30[15], temp29[15], temp28[15], temp27[15], temp26[15], temp25[15], temp24[15], temp23[15], temp22[15], temp21[15], temp20[15], temp19[15], temp18[15], temp17[15], temp16[15], temp15[15], temp14[15], temp13[15], temp12[15], temp11[15], temp10[15], temp9[15], temp8[15], temp7[15], temp6[15], temp5[15], temp4[15], temp3[15], temp2[15], temp1[15], temp0[15]}, in2[4:0], out[15]);
mux32to1 m16({temp31[16], temp30[16], temp29[16], temp28[16], temp27[16], temp26[16], temp25[16], temp24[16], temp23[16], temp22[16], temp21[16], temp20[16], temp19[16], temp18[16], temp17[16], temp16[16], temp15[16], temp14[16], temp13[16], temp12[16], temp11[16], temp10[16], temp9[16], temp8[16], temp7[16], temp6[16], temp5[16], temp4[16], temp3[16], temp2[16], temp1[16], temp0[16]}, in2[4:0], out[16]);
mux32to1 m17({temp31[17], temp30[17], temp29[17], temp28[17], temp27[17], temp26[17], temp25[17], temp24[17], temp23[17], temp22[17], temp21[17], temp20[17], temp19[17], temp18[17], temp17[17], temp16[17], temp15[17], temp14[17], temp13[17], temp12[17], temp11[17], temp10[17], temp9[17], temp8[17], temp7[17], temp6[17], temp5[17], temp4[17], temp3[17], temp2[17], temp1[17], temp0[17]}, in2[4:0], out[17]);
mux32to1 m18({temp31[18], temp30[18], temp29[18], temp28[18], temp27[18], temp26[18], temp25[18], temp24[18], temp23[18], temp22[18], temp21[18], temp20[18], temp19[18], temp18[18], temp17[18], temp16[18], temp15[18], temp14[18], temp13[18], temp12[18], temp11[18], temp10[18], temp9[18], temp8[18], temp7[18], temp6[18], temp5[18], temp4[18], temp3[18], temp2[18], temp1[18], temp0[18]}, in2[4:0], out[18]);
mux32to1 m19({temp31[19], temp30[19], temp29[19], temp28[19], temp27[19], temp26[19], temp25[19], temp24[19], temp23[19], temp22[19], temp21[19], temp20[19], temp19[19], temp18[19], temp17[19], temp16[19], temp15[19], temp14[19], temp13[19], temp12[19], temp11[19], temp10[19], temp9[19], temp8[19], temp7[19], temp6[19], temp5[19], temp4[19], temp3[19], temp2[19], temp1[19], temp0[19]}, in2[4:0], out[19]);
mux32to1 m20({temp31[20], temp30[20], temp29[20], temp28[20], temp27[20], temp26[20], temp25[20], temp24[20], temp23[20], temp22[20], temp21[20], temp20[20], temp19[20], temp18[20], temp17[20], temp16[20], temp15[20], temp14[20], temp13[20], temp12[20], temp11[20], temp10[20], temp9[20], temp8[20], temp7[20], temp6[20], temp5[20], temp4[20], temp3[20], temp2[20], temp1[20], temp0[20]}, in2[4:0], out[20]);
mux32to1 m21({temp31[21], temp30[21], temp29[21], temp28[21], temp27[21], temp26[21], temp25[21], temp24[21], temp23[21], temp22[21], temp21[21], temp20[21], temp19[21], temp18[21], temp17[21], temp16[21], temp15[21], temp14[21], temp13[21], temp12[21], temp11[21], temp10[21], temp9[21], temp8[21], temp7[21], temp6[21], temp5[21], temp4[21], temp3[21], temp2[21], temp1[21], temp0[21]}, in2[4:0], out[21]);
mux32to1 m22({temp31[22], temp30[22], temp29[22], temp28[22], temp27[22], temp26[22], temp25[22], temp24[22], temp23[22], temp22[22], temp21[22], temp20[22], temp19[22], temp18[22], temp17[22], temp16[22], temp15[22], temp14[22], temp13[22], temp12[22], temp11[22], temp10[22], temp9[22], temp8[22], temp7[22], temp6[22], temp5[22], temp4[22], temp3[22], temp2[22], temp1[22], temp0[22]}, in2[4:0], out[22]);
mux32to1 m23({temp31[23], temp30[23], temp29[23], temp28[23], temp27[23], temp26[23], temp25[23], temp24[23], temp23[23], temp22[23], temp21[23], temp20[23], temp19[23], temp18[23], temp17[23], temp16[23], temp15[23], temp14[23], temp13[23], temp12[23], temp11[23], temp10[23], temp9[23], temp8[23], temp7[23], temp6[23], temp5[23], temp4[23], temp3[23], temp2[23], temp1[23], temp0[23]}, in2[4:0], out[23]);
mux32to1 m24({temp31[24], temp30[24], temp29[24], temp28[24], temp27[24], temp26[24], temp25[24], temp24[24], temp23[24], temp22[24], temp21[24], temp20[24], temp19[24], temp18[24], temp17[24], temp16[24], temp15[24], temp14[24], temp13[24], temp12[24], temp11[24], temp10[24], temp9[24], temp8[24], temp7[24], temp6[24], temp5[24], temp4[24], temp3[24], temp2[24], temp1[24], temp0[24]}, in2[4:0], out[24]);
mux32to1 m25({temp31[25], temp30[25], temp29[25], temp28[25], temp27[25], temp26[25], temp25[25], temp24[25], temp23[25], temp22[25], temp21[25], temp20[25], temp19[25], temp18[25], temp17[25], temp16[25], temp15[25], temp14[25], temp13[25], temp12[25], temp11[25], temp10[25], temp9[25], temp8[25], temp7[25], temp6[25], temp5[25], temp4[25], temp3[25], temp2[25], temp1[25], temp0[25]}, in2[4:0], out[25]);
mux32to1 m26({temp31[26], temp30[26], temp29[26], temp28[26], temp27[26], temp26[26], temp25[26], temp24[26], temp23[26], temp22[26], temp21[26], temp20[26], temp19[26], temp18[26], temp17[26], temp16[26], temp15[26], temp14[26], temp13[26], temp12[26], temp11[26], temp10[26], temp9[26], temp8[26], temp7[26], temp6[26], temp5[26], temp4[26], temp3[26], temp2[26], temp1[26], temp0[26]}, in2[4:0], out[26]);
mux32to1 m27({temp31[27], temp30[27], temp29[27], temp28[27], temp27[27], temp26[27], temp25[27], temp24[27], temp23[27], temp22[27], temp21[27], temp20[27], temp19[27], temp18[27], temp17[27], temp16[27], temp15[27], temp14[27], temp13[27], temp12[27], temp11[27], temp10[27], temp9[27], temp8[27], temp7[27], temp6[27], temp5[27], temp4[27], temp3[27], temp2[27], temp1[27], temp0[27]}, in2[4:0], out[27]);
mux32to1 m28({temp31[28], temp30[28], temp29[28], temp28[28], temp27[28], temp26[28], temp25[28], temp24[28], temp23[28], temp22[28], temp21[28], temp20[28], temp19[28], temp18[28], temp17[28], temp16[28], temp15[28], temp14[28], temp13[28], temp12[28], temp11[28], temp10[28], temp9[28], temp8[28], temp7[28], temp6[28], temp5[28], temp4[28], temp3[28], temp2[28], temp1[28], temp0[28]}, in2[4:0], out[28]);
mux32to1 m29({temp31[29], temp30[29], temp29[29], temp28[29], temp27[29], temp26[29], temp25[29], temp24[29], temp23[29], temp22[29], temp21[29], temp20[29], temp19[29], temp18[29], temp17[29], temp16[29], temp15[29], temp14[29], temp13[29], temp12[29], temp11[29], temp10[29], temp9[29], temp8[29], temp7[29], temp6[29], temp5[29], temp4[29], temp3[29], temp2[29], temp1[29], temp0[29]}, in2[4:0], out[29]);
mux32to1 m30({temp31[30], temp30[30], temp29[30], temp28[30], temp27[30], temp26[30], temp25[30], temp24[30], temp23[30], temp22[30], temp21[30], temp20[30], temp19[30], temp18[30], temp17[30], temp16[30], temp15[30], temp14[30], temp13[30], temp12[30], temp11[30], temp10[30], temp9[30], temp8[30], temp7[30], temp6[30], temp5[30], temp4[30], temp3[30], temp2[30], temp1[30], temp0[30]}, in2[4:0], out[30]);
mux32to1 m31({temp31[31], temp30[31], temp29[31], temp28[31], temp27[31], temp26[31], temp25[31], temp24[31], temp23[31], temp22[31], temp21[31], temp20[31], temp19[31], temp18[31], temp17[31], temp16[31], temp15[31], temp14[31], temp13[31], temp12[31], temp11[31], temp10[31], temp9[31], temp8[31], temp7[31], temp6[31], temp5[31], temp4[31], temp3[31], temp2[31], temp1[31], temp0[31]}, in2[4:0], out[31]);

	 
	
endmodule